`timescale 1ns/10ps
module CLE ( clk, reset, rom_q, rom_a, sram_q, sram_a, sram_d, sram_wen, finish);
input         clk;
input         reset;
input  [7:0]  rom_q;
output [6:0]  rom_a;
input  [7:0]  sram_q;
output [9:0]  sram_a;
output [7:0]  sram_d;
output        sram_wen;
output        finish;

//parameter declaration
parameter IDLE      =2'd0;
parameter READ      =2'd1;
parameter PROCCESS  =2'd2;
parameter DONE      =2'd3;

//reg declaration

reg [6:0]   rom_a,    n_rom_a;
reg [9:0]   sram_a,   n_sram_a;
reg [7:0]   sram_d,   n_sram_d;
reg [1:0]   state,    next_state;
reg         sram_wen, n_sram_wen;
reg         finish,   n_finish;
reg         temp[0:1024];
reg [7:0]   count,n_count;
//combinational part
always@(*) begin
    n_finish = finish;
    n_count = count;
    n_sram_wen = sram_wen;
    n_sram_d = sram_d;
    n_sram_a = sram_a;
    n_rom_a = rom_a;
    case(state)
        IDLE: begin
            next_state = READ;
            n_rom_a = 0;
        end
        READ: begin   //iteration 128 times to read
            if(count < 128)begin
                for(i=0;i<8;i=i+1)
                    temp[8*count+i] = rom_q[i];
                n_count = count +1;
                n_rom_a = rom_a+1;
                next_state = READ;
            end
            else begin
                next_state = PROCESS;
        
            end
        end
        
        PROCCESS: begin
        end

        DONE: begin
        end

end

//sequential part
always@(posedge clk or posedge reset) begin
    if(reset) begin
        state <= IDLE;
        rom_a <= 0;
        sram_a <= 0;
        sram_d <= 0;
        sram_wen <= 0 ;
        finish <= 0;
        count <= 0
    end
    else begin
        state <= next_state;
        rom_a <= n_rom_a;
        sram_a <=n_sram_a;
        sram_d <=n_sram_d;
        sram_wem <=n_sram_wen;
        count <= n_count;
        finish <= n_finish;
    end
end
endmodule
